`ifndef _UDP_DEFINES_
 `define _UDP_DEFINES_ 1
 /**********************************************************
  * To add a register, 4 things need to be specified:
  * 1- block size, and block address
  * 2- Internal addresses used by the module internally
  * 3- External addresses to be used by test scripts
  * 4- Add the regs to the display command to easily get addresses
  * 
  * please see NF_2.1_defines.v for an example
  **********************************************************/

 /**********************************************************
  * The UDP address space is divided into classes:
  *      - 4096 blocks of size 64 words
  *      - 256  blocks of size 1k words
  * FIXME: Any addresses that begin with 3 zeros are size 32 blocks
  * FIXME: All other addresses belong to blocks of size 512
  **********************************************************/

 // --- Define address ranges
 // 12 bits to identify blocks of size 64
 `define UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH  12
 `define UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH    6
 `define UDP_BLOCK_SIZE_64_TAG               ({(`UDP_REG_ADDR_WIDTH-`UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH-`UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH){1'b0}})

 // 8 bits to identify blocks of size 1k words
 `define UDP_BLOCK_SIZE_1k_BLOCK_ADDR_WIDTH   8
 `define UDP_BLOCK_SIZE_1k_REG_ADDR_WIDTH     10
 `define UDP_BLOCK_SIZE_1k_TAG               ({{(`UDP_REG_ADDR_WIDTH-`UDP_BLOCK_SIZE_1k_BLOCK_ADDR_WIDTH-`UDP_BLOCK_SIZE_1k_REG_ADDR_WIDTH-1){1'b0}}, 1'b1})

 // --- Define subblock address ranges
 //
 // These are splits of the 64 address range
 `define UDP_SUB_BLOCK_SIZE_32_BLOCK_ADDR_WIDTH  1
 `define UDP_SUB_BLOCK_SIZE_32_REG_ADDR_WIDTH    5

 // --- Size 64 Block register addresses
 `define OP_LUT_REG_ADDR_WIDTH           `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define OP_LUT_BLOCK_ADDR_WIDTH         `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define OP_LUT_BLOCK_ADDR               `OP_LUT_BLOCK_ADDR_WIDTH'h1
 `define OP_LUT_BLOCK_TAG                ({`UDP_BLOCK_SIZE_64_TAG, `OP_LUT_BLOCK_ADDR})

 `define OP_LUT_NON_CNTR_REG_ADDR_WIDTH    `UDP_SUB_BLOCK_SIZE_32_REG_ADDR_WIDTH
 `define OP_LUT_NON_CNTR_BLOCK_ADDR_WIDTH  `UDP_SUB_BLOCK_SIZE_32_BLOCK_ADDR_WIDTH
 `define OP_LUT_NON_CNTR_BLOCK_ADDR        `OP_LUT_NON_CNTR_BLOCK_ADDR_WIDTH'h0
 `define OP_LUT_NON_CNTR_BLOCK_TAG         ({`OP_LUT_BLOCK_TAG, `OP_LUT_NON_CNTR_BLOCK_ADDR})

 `define OP_LUT_CNTR_REG_ADDR_WIDTH        `UDP_SUB_BLOCK_SIZE_32_REG_ADDR_WIDTH
 `define OP_LUT_CNTR_BLOCK_ADDR_WIDTH      `UDP_SUB_BLOCK_SIZE_32_BLOCK_ADDR_WIDTH
 `define OP_LUT_CNTR_BLOCK_ADDR            `OP_LUT_CNTR_BLOCK_ADDR_WIDTH'h1
 `define OP_LUT_CNTR_BLOCK_TAG             ({`OP_LUT_BLOCK_TAG, `OP_LUT_CNTR_BLOCK_ADDR})

 `define IN_ARB_REG_ADDR_WIDTH           `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define IN_ARB_BLOCK_ADDR_WIDTH         `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define IN_ARB_BLOCK_ADDR               `IN_ARB_BLOCK_ADDR_WIDTH'h2
 `define IN_ARB_BLOCK_TAG                ({`UDP_BLOCK_SIZE_64_TAG, `IN_ARB_BLOCK_ADDR})

 `define EVT_CAP_REG_ADDR_WIDTH          `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define EVT_CAP_BLOCK_ADDR_WIDTH        `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define EVT_CAP_BLOCK_ADDR              `EVT_CAP_BLOCK_ADDR_WIDTH'h3
 `define EVT_CAP_BLOCK_TAG               ({`UDP_BLOCK_SIZE_64_TAG, `EVT_CAP_BLOCK_ADDR})

 `define RATE_LIMIT_REG_ADDR_WIDTH       `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define RATE_LIMIT_BLOCK_ADDR_WIDTH     `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define RATE_LIMIT_BLOCK_ADDR           `RATE_LIMIT_BLOCK_ADDR_WIDTH'h4
 `define RATE_LIMIT_BLOCK_TAG            ({`UDP_BLOCK_SIZE_64_TAG, `RATE_LIMIT_BLOCK_ADDR})

 `define DELAY_REG_ADDR_WIDTH            `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define DELAY_BLOCK_ADDR_WIDTH          `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define DELAY_BLOCK_ADDR                `DELAY_BLOCK_ADDR_WIDTH'h5
 `define DELAY_BLOCK_TAG                 ({`UDP_BLOCK_SIZE_64_TAG, `DELAY_BLOCK_ADDR})

 `define SWITCH_OP_LUT_REG_ADDR_WIDTH    `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define SWITCH_OP_LUT_BLOCK_ADDR_WIDTH  `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define SWITCH_OP_LUT_BLOCK_ADDR        `SWITCH_OP_LUT_BLOCK_ADDR_WIDTH'h6
 `define SWITCH_OP_LUT_BLOCK_TAG         ({`UDP_BLOCK_SIZE_64_TAG, `SWITCH_OP_LUT_BLOCK_ADDR})

 `define BRAM_OQ_REG_ADDR_WIDTH          `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define BRAM_OQ_BLOCK_ADDR_WIDTH        `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define BRAM_OQ_BLOCK_ADDR              `BRAM_OQ_BLOCK_ADDR_WIDTH'h7
 `define BRAM_OQ_BLOCK_TAG               ({`UDP_BLOCK_SIZE_64_TAG, `BRAM_OQ_BLOCK_ADDR})

 `define RCP_REG_ADDR_WIDTH               `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define RCP_BLOCK_ADDR_WIDTH             `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define RCP_BLOCK_ADDR                   `RCP_BLOCK_ADDR_WIDTH'h8
 `define RCP_BLOCK_TAG                    ({`UDP_BLOCK_SIZE_64_TAG, `RCP_BLOCK_ADDR})


 `define ENCAP_REG_ADDR_WIDTH               `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define ENCAP_BLOCK_ADDR_WIDTH             `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define ENCAP_BLOCK_ADDR                   `RCP_BLOCK_ADDR_WIDTH'h9
 `define ENCAP_BLOCK_TAG                    ({`UDP_BLOCK_SIZE_64_TAG, `ENCAP_BLOCK_ADDR})

 `define DECAP_REG_ADDR_WIDTH               `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define DECAP_BLOCK_ADDR_WIDTH             `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define DECAP_BLOCK_ADDR                   `RCP_BLOCK_ADDR_WIDTH'hA
 `define DECAP_BLOCK_TAG                    ({`UDP_BLOCK_SIZE_64_TAG, `DECAP_BLOCK_ADDR})



 `define PKT_GEN_CTRL_REG_ADDR_WIDTH     `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define PKT_GEN_CTRL_BLOCK_ADDR_WIDTH   `UDP_BLOCK_SIZE_64_BLOCK_ADDR_WIDTH
 `define PKT_GEN_CTRL_BLOCK_ADDR         `EVT_CAP_BLOCK_ADDR_WIDTH'hB
 `define PKT_GEN_CTRL_BLOCK_TAG          ({`UDP_BLOCK_SIZE_64_TAG, `EVT_CAP_BLOCK_ADDR})


 // --- Size 1024 Block register addresses
 `define OQ_REG_ADDR_WIDTH               `UDP_BLOCK_SIZE_1k_REG_ADDR_WIDTH
 `define OQ_BLOCK_ADDR_WIDTH             `UDP_BLOCK_SIZE_1k_BLOCK_ADDR_WIDTH
 `define OQ_BLOCK_ADDR                   `OQ_BLOCK_ADDR_WIDTH'h1
 `define OQ_BLOCK_TAG                    ({`UDP_BLOCK_SIZE_1k_TAG, `OQ_BLOCK_ADDR})



 // 1- add additional blocks here



 /*******************************************************************
  -- Internal addresses -- these are used inside the modules
  *******************************************************************/
 // --- inut arbiter internal regs
 `define IN_ARB_NUM_PKTS_SENT            `IN_ARB_REG_ADDR_WIDTH'h0
 `define IN_ARB_LAST_PKT_WORD_0_LO       `IN_ARB_REG_ADDR_WIDTH'h1
 `define IN_ARB_LAST_PKT_WORD_0_HI       `IN_ARB_REG_ADDR_WIDTH'h2
 `define IN_ARB_LAST_PKT_CTRL_0          `IN_ARB_REG_ADDR_WIDTH'h3
 `define IN_ARB_LAST_PKT_WORD_1_LO       `IN_ARB_REG_ADDR_WIDTH'h4
 `define IN_ARB_LAST_PKT_WORD_1_HI       `IN_ARB_REG_ADDR_WIDTH'h5
 `define IN_ARB_LAST_PKT_CTRL_1          `IN_ARB_REG_ADDR_WIDTH'h6
 `define IN_ARB_STATE                    `IN_ARB_REG_ADDR_WIDTH'h7

 // --- switch output port lut internal reg addresses
 `define SWITCH_OP_LUT_PORTS_MAC_HI      `SWITCH_OP_LUT_REG_ADDR_WIDTH'h0
 `define SWITCH_OP_LUT_MAC_LO            `SWITCH_OP_LUT_REG_ADDR_WIDTH'h1
 `define SWITCH_OP_LUT_NUM_HITS          `SWITCH_OP_LUT_REG_ADDR_WIDTH'h2
 `define SWITCH_OP_LUT_NUM_MISSES        `SWITCH_OP_LUT_REG_ADDR_WIDTH'h3
 `define SWITCH_OP_LUT_MAC_LUT_RD_ADDR   `SWITCH_OP_LUT_REG_ADDR_WIDTH'h4
 `define SWITCH_OP_LUT_MAC_LUT_WR_ADDR   `SWITCH_OP_LUT_REG_ADDR_WIDTH'h5

 // --- router output port lut internal reg addresses
 /* Define table sizes */
 `define ROUTER_RT_SIZE                  32
 `define ROUTER_ARP_SIZE                 32
 `define ROUTER_DST_IP_FILTER_TABLE_DEPTH 32

 /* Access to the ARP table */
 `define ROUTER_OP_LUT_ARP_MAC_HI        `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h0
 `define ROUTER_OP_LUT_ARP_MAC_LO        `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h1
 `define ROUTER_OP_LUT_ARP_NEXT_HOP_IP   `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h2
 `define ROUTER_OP_LUT_ARP_LUT_RD_ADDR   `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h3
 `define ROUTER_OP_LUT_ARP_LUT_WR_ADDR   `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h4

 /* Access to the Routing Table */
 `define ROUTER_OP_LUT_RT_IP             `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h5
 `define ROUTER_OP_LUT_RT_MASK           `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h6
 `define ROUTER_OP_LUT_RT_NEXT_HOP_IP    `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h7
 `define ROUTER_OP_LUT_RT_OUTPUT_PORT    `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h8
 `define ROUTER_OP_LUT_RT_LUT_RD_ADDR    `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h9
 `define ROUTER_OP_LUT_RT_LUT_WR_ADDR    `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'ha

 /* Stats counters */
 `define ROUTER_OP_LUT_ARP_NUM_MISSES    `OP_LUT_CNTR_REG_ADDR_WIDTH'h0
 `define ROUTER_OP_LUT_LPM_NUM_MISSES    `OP_LUT_CNTR_REG_ADDR_WIDTH'h1
 `define ROUTER_OP_LUT_NUM_CPU_PKTS_SENT `OP_LUT_CNTR_REG_ADDR_WIDTH'h2
 `define ROUTER_OP_LUT_NUM_BAD_OPTS_VER  `OP_LUT_CNTR_REG_ADDR_WIDTH'h3
 `define ROUTER_OP_LUT_NUM_BAD_CHKSUMS   `OP_LUT_CNTR_REG_ADDR_WIDTH'h4
 `define ROUTER_OP_LUT_NUM_BAD_TTLS      `OP_LUT_CNTR_REG_ADDR_WIDTH'h5
 `define ROUTER_OP_LUT_NUM_NON_IP_RCVD   `OP_LUT_CNTR_REG_ADDR_WIDTH'h6
 `define ROUTER_OP_LUT_NUM_PKTS_FORWARDED `OP_LUT_CNTR_REG_ADDR_WIDTH'h7
 `define ROUTER_OP_LUT_NUM_WRONG_DEST    `OP_LUT_CNTR_REG_ADDR_WIDTH'h8
 `define ROUTER_OP_LUT_NUM_FILTERED_PKTS `OP_LUT_CNTR_REG_ADDR_WIDTH'h9

 /*ENCAP Module */
 `define ENCAP_ENABLE                      `ENCAP_REG_ADDR_WIDTH'h2
 `define ENCAP_IP_DATA_0                   `ENCAP_REG_ADDR_WIDTH'h3
 `define ENCAP_IP_DATA_1                   `ENCAP_REG_ADDR_WIDTH'h4
 `define ENCAP_IP_DATA_2                   `ENCAP_REG_ADDR_WIDTH'h5
 `define ENCAP_IP_DATA_3                   `ENCAP_REG_ADDR_WIDTH'h6
 `define ENCAP_IP_DATA_4                   `ENCAP_REG_ADDR_WIDTH'h7
 `define ENCAP_IP_DATA_5                   `ENCAP_REG_ADDR_WIDTH'h8
 `define ENCAP_NUM_PACKET_IN               `ENCAP_REG_ADDR_WIDTH'h9
 `define ENCAP_NUM_PACKET_OUT              `ENCAP_REG_ADDR_WIDTH'ha
 `define ENCAP_NUM_BYTES_IN                `ENCAP_REG_ADDR_WIDTH'hb
 `define ENCAP_NUM_BYTES_OUT               `ENCAP_REG_ADDR_WIDTH'hc

 /*DECAP Module */
 `define DECAP_NUM_WORD_IN                  `DECAP_REG_ADDR_WIDTH'h4
 `define DECAP_NUM_WORD_OUT                 `DECAP_REG_ADDR_WIDTH'h5
 `define DECAP_VALID_TUNNELING              `DECAP_REG_ADDR_WIDTH'h6
 `define DECAP_USER_DATA_PATH_HEADER        `DECAP_REG_ADDR_WIDTH'h7
 `define DECAP_NUM_PACKET_IN                `DECAP_REG_ADDR_WIDTH'h8
 `define DECAP_NUM_PACKET_OUT               `DECAP_REG_ADDR_WIDTH'h9



 /* Config registers */
 // high 16 bits of MAC address of MAC port 0
 `define ROUTER_OP_LUT_MAC_0_HI          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'hb
 // low 32 bits of MAC address of MAC port 0
 `define ROUTER_OP_LUT_MAC_0_LO          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'hc

 // high 16 bits of MAC address of MAC port 1
 `define ROUTER_OP_LUT_MAC_1_HI          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'hd
 // low 32 bits of MAC address of MAC port 1
 `define ROUTER_OP_LUT_MAC_1_LO          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'he

 // high 16 bits of MAC address of MAC port 2
 `define ROUTER_OP_LUT_MAC_2_HI          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'hf
 // low 32 bits of MAC address of MAC port 2
 `define ROUTER_OP_LUT_MAC_2_LO          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h10

 // high 16 bits of MAC address of MAC port 3
 `define ROUTER_OP_LUT_MAC_3_HI          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h11
 // low 32 bits of MAC address of MAC port 3
 `define ROUTER_OP_LUT_MAC_3_LO          `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h12

 /* Access to the destination ip filter */
 `define ROUTER_OP_LUT_DST_IP_FILTER_IP      `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h13
 `define ROUTER_OP_LUT_DST_IP_FILTER_RD_ADDR `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h14
 `define ROUTER_OP_LUT_DST_IP_FILTER_WR_ADDR `OP_LUT_NON_CNTR_REG_ADDR_WIDTH'h15

 `define DEFAULT_MAC_0_HI                32'h0000_cafe
 `define DEFAULT_MAC_0_LO                32'hf00d_0001
 `define DEFAULT_MAC_1_HI                32'h0000_cafe
 `define DEFAULT_MAC_1_LO                32'hf00d_0002
 `define DEFAULT_MAC_2_HI                32'h0000_cafe
 `define DEFAULT_MAC_2_LO                32'hf00d_0003
 `define DEFAULT_MAC_3_HI                32'h0000_cafe
 `define DEFAULT_MAC_3_LO                32'hf00d_0004

 // --- output queues internal registers
 // 
 // Note: OQ_REG_HELPER_BLOCK_ADDR_WIDTH must be calculated manually... sigh
 `define OQ_REG_HELPER_ADDR_WIDTH        `UDP_BLOCK_SIZE_64_REG_ADDR_WIDTH
 `define OQ_REG_HELPER_BLOCK_ADDR_WIDTH  4

 `define OQ_NUM_WORDS_LEFT               `OQ_REG_HELPER_ADDR_WIDTH'h0
 `define OQ_NUM_PKT_BYTES_STORED         `OQ_REG_HELPER_ADDR_WIDTH'h1
 `define OQ_NUM_OVERHEAD_BYTES_STORED    `OQ_REG_HELPER_ADDR_WIDTH'h2
 `define OQ_NUM_PKTS_STORED              `OQ_REG_HELPER_ADDR_WIDTH'h3
 `define OQ_NUM_PKTS_DROPPED             `OQ_REG_HELPER_ADDR_WIDTH'h4
 `define OQ_NUM_PKT_BYTES_REMOVED        `OQ_REG_HELPER_ADDR_WIDTH'h5
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED   `OQ_REG_HELPER_ADDR_WIDTH'h6
 `define OQ_NUM_PKTS_REMOVED             `OQ_REG_HELPER_ADDR_WIDTH'h7
 `define OQ_ADDRESS_HI                   `OQ_REG_HELPER_ADDR_WIDTH'h8
 `define OQ_ADDRESS_LO                   `OQ_REG_HELPER_ADDR_WIDTH'h9
 `define OQ_WR_ADDRESS                   `OQ_REG_HELPER_ADDR_WIDTH'ha
 `define OQ_RD_ADDRESS                   `OQ_REG_HELPER_ADDR_WIDTH'hb
 `define OQ_NUM_PKTS_IN_Q                `OQ_REG_HELPER_ADDR_WIDTH'hc
 `define OQ_MAX_PKTS_IN_Q                `OQ_REG_HELPER_ADDR_WIDTH'hd
 `define OQ_CONTROL                      `OQ_REG_HELPER_ADDR_WIDTH'he
 `define OQ_NUM_WORDS_IN_Q               `OQ_REG_HELPER_ADDR_WIDTH'hf
 `define OQ_FULL_THRESH                  `OQ_REG_HELPER_ADDR_WIDTH'h10
 ////////////////////////////////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT                `OQ_REG_HELPER_ADDR_WIDTH'h11
 `define JAN_OQ_PKTRM_CNT                `OQ_REG_HELPER_ADDR_WIDTH'h12
 `define JAN_OQ_AB_STATE                 `OQ_REG_HELPER_ADDR_WIDTH'h13
 `define JAN_OQ_AB_MOD_STATE             `OQ_REG_HELPER_ADDR_WIDTH'h14
 `define JAN_OQ_AC_STATE                 `OQ_REG_HELPER_ADDR_WIDTH'h15
 `define JAN_OQ_AC_MOD_STATE             `OQ_REG_HELPER_ADDR_WIDTH'h16

///////////////////////////////////////////////////////////////////////////////
 // Each SRAM is 2MB (512k x 36 bits)
 // Carve it up to equal parts for each output queue
 `define OQ_DEFAULT_ADDR_LOW(j, num_oqs)  ((j)*20'h8_0000/(num_oqs))
 `define OQ_DEFAULT_ADDR_HIGH(j, num_oqs) (((j+1)*20'h8_0000/(num_oqs)) - 1)

 `define OQ_DEFAULT_MAX_PKTS              32'hffff_ffff

 `define OQ_ENABLE_SEND_BIT              `OP_LUT_REG_ADDR_WIDTH'h1
 `define OQ_INITIALIZE_OQ_BIT            `OP_LUT_REG_ADDR_WIDTH'h2
 `define OQ_ENABLE_SEND_BIT_NUM          0
 `define OQ_INITIALIZE_OQ_BIT_NUM        1

 // --- Delay registers
 `define DELAY_ENABLE                    `DELAY_REG_ADDR_WIDTH'h0
 `define DELAY_LENGTH                    `DELAY_REG_ADDR_WIDTH'h1
 `define DELAY_1ST_WORD_HI               `DELAY_REG_ADDR_WIDTH'h2
 `define DELAY_1ST_WORD_LO               `DELAY_REG_ADDR_WIDTH'h3


 // --- Rate limiter registers
 `define RATE_LIMIT_ENABLE               `RATE_LIMIT_REG_ADDR_WIDTH'h0
 `define RATE_LIMIT_SHIFT                `RATE_LIMIT_REG_ADDR_WIDTH'h1

 // --- event capture internal regs
 `define EVT_CAP_ENABLE_CAPTURE          `EVT_CAP_REG_ADDR_WIDTH'h0
 `define EVT_CAP_SEND_PKT                `EVT_CAP_REG_ADDR_WIDTH'h1
 `define EVT_CAP_DST_MAC_HI              `EVT_CAP_REG_ADDR_WIDTH'h2
 `define EVT_CAP_DST_MAC_LO              `EVT_CAP_REG_ADDR_WIDTH'h3
 `define EVT_CAP_SRC_MAC_HI              `EVT_CAP_REG_ADDR_WIDTH'h4
 `define EVT_CAP_SRC_MAC_LO              `EVT_CAP_REG_ADDR_WIDTH'h5
 `define EVT_CAP_ETHERTYPE               `EVT_CAP_REG_ADDR_WIDTH'h6
 `define EVT_CAP_IP_DST                  `EVT_CAP_REG_ADDR_WIDTH'h7
 `define EVT_CAP_IP_SRC                  `EVT_CAP_REG_ADDR_WIDTH'h8
 `define EVT_CAP_MONITOR_MASK            `EVT_CAP_REG_ADDR_WIDTH'h9
 `define EVT_CAP_SIGNAL_ID_MASK          `EVT_CAP_REG_ADDR_WIDTH'ha
 `define EVT_CAP_NUM_EVTS_DROPPED        `EVT_CAP_REG_ADDR_WIDTH'hb
 `define EVT_CAP_UDP_SRC_PORT            `EVT_CAP_REG_ADDR_WIDTH'hc
 `define EVT_CAP_UDP_DST_PORT            `EVT_CAP_REG_ADDR_WIDTH'hd
 `define EVT_CAP_OUTPUT_PORTS            `EVT_CAP_REG_ADDR_WIDTH'he
 `define EVT_CAP_RESET_TIMERS            `EVT_CAP_REG_ADDR_WIDTH'hf
 `define EVT_CAP_TIMER_RESOLUTION        `EVT_CAP_REG_ADDR_WIDTH'h10
 `define EVT_CAP_NUM_EVT_PKTS_SENT       `EVT_CAP_REG_ADDR_WIDTH'h11
 `define EVT_CAP_NUM_EVTS_SENT           `EVT_CAP_REG_ADDR_WIDTH'h12

 // --- Block RAM output queues
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_0  `BRAM_OQ_REG_ADDR_WIDTH'h0
 `define BRAM_OQ_NUM_PKTS_RECEIVED_0       `BRAM_OQ_REG_ADDR_WIDTH'h1
 `define BRAM_OQ_NUM_PKTS_DROPPED_0        `BRAM_OQ_REG_ADDR_WIDTH'h2
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_1  `BRAM_OQ_REG_ADDR_WIDTH'h3
 `define BRAM_OQ_NUM_PKTS_RECEIVED_1       `BRAM_OQ_REG_ADDR_WIDTH'h4
 `define BRAM_OQ_NUM_PKTS_DROPPED_1        `BRAM_OQ_REG_ADDR_WIDTH'h5
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_2  `BRAM_OQ_REG_ADDR_WIDTH'h6
 `define BRAM_OQ_NUM_PKTS_RECEIVED_2       `BRAM_OQ_REG_ADDR_WIDTH'h7
 `define BRAM_OQ_NUM_PKTS_DROPPED_2        `BRAM_OQ_REG_ADDR_WIDTH'h8
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_3  `BRAM_OQ_REG_ADDR_WIDTH'h9
 `define BRAM_OQ_NUM_PKTS_RECEIVED_3       `BRAM_OQ_REG_ADDR_WIDTH'ha
 `define BRAM_OQ_NUM_PKTS_DROPPED_3        `BRAM_OQ_REG_ADDR_WIDTH'hb
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_4  `BRAM_OQ_REG_ADDR_WIDTH'hc
 `define BRAM_OQ_NUM_PKTS_RECEIVED_4       `BRAM_OQ_REG_ADDR_WIDTH'hd
 `define BRAM_OQ_NUM_PKTS_DROPPED_4        `BRAM_OQ_REG_ADDR_WIDTH'he
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_5  `BRAM_OQ_REG_ADDR_WIDTH'hf
 `define BRAM_OQ_NUM_PKTS_RECEIVED_5       `BRAM_OQ_REG_ADDR_WIDTH'h10
 `define BRAM_OQ_NUM_PKTS_DROPPED_5        `BRAM_OQ_REG_ADDR_WIDTH'h11
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_6  `BRAM_OQ_REG_ADDR_WIDTH'h12
 `define BRAM_OQ_NUM_PKTS_RECEIVED_6       `BRAM_OQ_REG_ADDR_WIDTH'h13
 `define BRAM_OQ_NUM_PKTS_DROPPED_6        `BRAM_OQ_REG_ADDR_WIDTH'h14
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_7  `BRAM_OQ_REG_ADDR_WIDTH'h15
 `define BRAM_OQ_NUM_PKTS_RECEIVED_7       `BRAM_OQ_REG_ADDR_WIDTH'h16
 `define BRAM_OQ_NUM_PKTS_DROPPED_7        `BRAM_OQ_REG_ADDR_WIDTH'h17
 `define BRAM_OQ_DISABLE_QUEUES            `BRAM_OQ_REG_ADDR_WIDTH'h18
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_0      `BRAM_OQ_REG_ADDR_WIDTH'h19
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_1      `BRAM_OQ_REG_ADDR_WIDTH'h1a
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_2      `BRAM_OQ_REG_ADDR_WIDTH'h1b
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_3      `BRAM_OQ_REG_ADDR_WIDTH'h1c
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_4      `BRAM_OQ_REG_ADDR_WIDTH'h1d
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_5      `BRAM_OQ_REG_ADDR_WIDTH'h1e
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_6      `BRAM_OQ_REG_ADDR_WIDTH'h1f
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_7      `BRAM_OQ_REG_ADDR_WIDTH'h20
 
 //-- RCP registers
 `define RCP_RATE                        `RCP_REG_ADDR_WIDTH'h2
 `define RCP_MAC_0_RTT_L                 `RCP_REG_ADDR_WIDTH'h4
 `define RCP_MAC_0_RTT_H                 `RCP_REG_ADDR_WIDTH'h5
 `define RCP_MAC_0_NUM_RCP               `RCP_REG_ADDR_WIDTH'h6
 `define RCP_MAC_0_NUM_BYTE_L            `RCP_REG_ADDR_WIDTH'h7
 `define RCP_MAC_0_NUM_BYTE_H            `RCP_REG_ADDR_WIDTH'h8
 `define RCP_MAC_1_RTT_L                 `RCP_REG_ADDR_WIDTH'h9
 `define RCP_MAC_1_RTT_H                 `RCP_REG_ADDR_WIDTH'ha
 `define RCP_MAC_1_NUM_RCP               `RCP_REG_ADDR_WIDTH'hb
 `define RCP_MAC_1_NUM_BYTE_L            `RCP_REG_ADDR_WIDTH'hc
 `define RCP_MAC_1_NUM_BYTE_H            `RCP_REG_ADDR_WIDTH'hd
 `define RCP_MAC_2_RTT_L                 `RCP_REG_ADDR_WIDTH'he
 `define RCP_MAC_2_RTT_H                 `RCP_REG_ADDR_WIDTH'hf
 `define RCP_MAC_2_NUM_RCP               `RCP_REG_ADDR_WIDTH'h10
 `define RCP_MAC_2_NUM_BYTE_L            `RCP_REG_ADDR_WIDTH'h11
 `define RCP_MAC_2_NUM_BYTE_H            `RCP_REG_ADDR_WIDTH'h12
 `define RCP_MAC_3_RTT_L                 `RCP_REG_ADDR_WIDTH'h13
 `define RCP_MAC_3_RTT_H                 `RCP_REG_ADDR_WIDTH'h14
 `define RCP_MAC_3_NUM_RCP               `RCP_REG_ADDR_WIDTH'h15
 `define RCP_MAC_3_NUM_BYTE_L            `RCP_REG_ADDR_WIDTH'h16
 `define RCP_MAC_3_NUM_BYTE_H            `RCP_REG_ADDR_WIDTH'h17

 // 2- add other internal addresses here


 /************************
   --- External addresses
  ************************/

 `define IN_ARB_NUM_PKTS_SENT_REG             (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_NUM_PKTS_SENT})
 `define IN_ARB_LAST_PKT_WORD_0_LO_REG        (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_WORD_0_LO})
 `define IN_ARB_LAST_PKT_WORD_0_HI_REG        (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_WORD_0_HI})
 `define IN_ARB_LAST_PKT_CTRL_0_REG           (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_CTRL_0   })
 `define IN_ARB_LAST_PKT_WORD_1_LO_REG        (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_WORD_1_LO})
 `define IN_ARB_LAST_PKT_WORD_1_HI_REG        (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_WORD_1_HI})
 `define IN_ARB_LAST_PKT_CTRL_1_REG           (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_LAST_PKT_CTRL_1   })
 `define IN_ARB_STATE_REG                     (`UDP_BASE_ADDRESS | {`IN_ARB_BLOCK_TAG, `IN_ARB_STATE   })

 `define SWITCH_OP_LUT_PORTS_MAC_HI_REG       (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_PORTS_MAC_HI})
 `define SWITCH_OP_LUT_MAC_LO_REG             (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_MAC_LO})
 `define SWITCH_OP_LUT_NUM_HITS_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_NUM_HITS})
 `define SWITCH_OP_LUT_NUM_MISSES_REG         (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_NUM_MISSES})
 `define SWITCH_OP_LUT_MAC_LUT_RD_ADDR_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_MAC_LUT_RD_ADDR})
 `define SWITCH_OP_LUT_MAC_LUT_WR_ADDR_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_BLOCK_TAG, `SWITCH_OP_LUT_MAC_LUT_WR_ADDR})

 `define ROUTER_OP_LUT_ARP_MAC_HI_REG         (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_MAC_HI})
 `define ROUTER_OP_LUT_ARP_MAC_LO_REG         (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_MAC_LO})
 `define ROUTER_OP_LUT_ARP_NEXT_HOP_IP_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_NEXT_HOP_IP})
 `define ROUTER_OP_LUT_ARP_LUT_RD_ADDR_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_LUT_RD_ADDR})
 `define ROUTER_OP_LUT_ARP_LUT_WR_ADDR_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_LUT_WR_ADDR})
 `define ROUTER_OP_LUT_RT_IP_REG              (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_IP})
 `define ROUTER_OP_LUT_RT_MASK_REG            (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_MASK})
 `define ROUTER_OP_LUT_RT_NEXT_HOP_IP_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_NEXT_HOP_IP})
 `define ROUTER_OP_LUT_RT_OUTPUT_PORT_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_OUTPUT_PORT})
 `define ROUTER_OP_LUT_RT_LUT_RD_ADDR_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_LUT_RD_ADDR})
 `define ROUTER_OP_LUT_RT_LUT_WR_ADDR_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_RT_LUT_WR_ADDR})
 `define ROUTER_OP_LUT_MAC_0_HI_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_0_HI})
 `define ROUTER_OP_LUT_MAC_0_LO_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_0_LO})
 `define ROUTER_OP_LUT_MAC_1_HI_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_1_HI})
 `define ROUTER_OP_LUT_MAC_1_LO_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_1_LO})
 `define ROUTER_OP_LUT_MAC_2_HI_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_2_HI})
 `define ROUTER_OP_LUT_MAC_2_LO_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_2_LO})
 `define ROUTER_OP_LUT_MAC_3_HI_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_3_HI})
 `define ROUTER_OP_LUT_MAC_3_LO_REG           (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_MAC_3_LO})
 `define ROUTER_OP_LUT_DST_IP_FILTER_IP_REG   (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_DST_IP_FILTER_IP})
 `define ROUTER_OP_LUT_DST_IP_FILTER_RD_ADDR_REG (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_DST_IP_FILTER_RD_ADDR})
 `define ROUTER_OP_LUT_DST_IP_FILTER_WR_ADDR_REG (`UDP_BASE_ADDRESS | {`OP_LUT_NON_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_DST_IP_FILTER_WR_ADDR})

 `define ROUTER_OP_LUT_ARP_NUM_MISSES_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_ARP_NUM_MISSES})
 `define ROUTER_OP_LUT_LPM_NUM_MISSES_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_LPM_NUM_MISSES})
 `define ROUTER_OP_LUT_NUM_CPU_PKTS_SENT_REG  (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_CPU_PKTS_SENT})
 `define ROUTER_OP_LUT_NUM_BAD_OPTS_VER_REG   (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_BAD_OPTS_VER})
 `define ROUTER_OP_LUT_NUM_BAD_CHKSUMS_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_BAD_CHKSUMS})
 `define ROUTER_OP_LUT_NUM_BAD_TTLS_REG       (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_BAD_TTLS})
 `define ROUTER_OP_LUT_NUM_NON_IP_RCVD_REG    (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_NON_IP_RCVD})
 `define ROUTER_OP_LUT_NUM_PKTS_FORWARDED_REG (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_PKTS_FORWARDED})
 `define ROUTER_OP_LUT_NUM_WRONG_DEST_REG     (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_WRONG_DEST})
 `define ROUTER_OP_LUT_NUM_FILTERED_PKTS_REG  (`UDP_BASE_ADDRESS | {`OP_LUT_CNTR_BLOCK_TAG, `ROUTER_OP_LUT_NUM_FILTERED_PKTS})

 `define OQ_NUM_WORDS_LEFT_REG_0              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_0        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_0   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_0             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_0            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_0       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_0  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_0            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_0                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_0                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_0                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_0                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_0               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_0               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_0                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_0                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_0              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG0                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG0                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG0                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG0             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG0                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG0             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_1              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_1        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_1   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_1             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_1            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_1       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_1  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_1            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_1                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_1                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_1                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_1                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_1               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_1               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_1                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_1                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_1              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h1}, `OQ_NUM_WORDS_IN_Q})
   //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG1                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG1                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG1                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG1             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG1                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_2              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_2        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_2   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_2             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_2            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_2       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_2  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_2            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_2                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_2                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_2                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_2                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_2               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_2               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_2                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_2                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_2              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h2}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG2                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG2                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG2                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG2             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG2                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG2             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_3              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_3        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_3   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_3             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_3            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_3       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_3  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_3            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_3                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_3                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_3                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_3                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_3               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_3               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_3                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_3                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_3              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h3}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG3                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG3                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG3                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG3             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG3                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG3             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_4              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_4        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_4   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_4             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_4            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_4       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_4  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_4            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_4                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_4                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_4                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_4                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_4               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_4               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_4                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_4                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_4              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h4}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG4                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG4                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG4                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG4             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG4                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG4             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_5              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_5        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_5   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_5             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_5            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_5       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_5  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_5            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_5                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_5                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_5                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_5                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_5               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_5               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_5                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_5                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_5              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h5}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG5                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG5                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG5                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG5             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG5                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG5             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////
 
 `define OQ_NUM_WORDS_LEFT_REG_6              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_6        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_6   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_6             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_6            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_6       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_6  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_6            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_6                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_6                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_6                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_6                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_6               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_6               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_6                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_6                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_6              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h6}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG6                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG6                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG6                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG6             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG6                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG6             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define OQ_NUM_WORDS_LEFT_REG_7              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_WORDS_LEFT})
 `define OQ_NUM_PKT_BYTES_STORED_REG_7        (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKT_BYTES_STORED})
 `define OQ_NUM_OVERHEAD_BYTES_STORED_REG_7   (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_OVERHEAD_BYTES_STORED})
 `define OQ_NUM_PKTS_STORED_REG_7             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKTS_STORED})
 `define OQ_NUM_PKTS_DROPPED_REG_7            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKTS_DROPPED})
 `define OQ_NUM_PKT_BYTES_REMOVED_REG_7       (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKT_BYTES_REMOVED})
 `define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_7  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_OVERHEAD_BYTES_REMOVED})
 `define OQ_NUM_PKTS_REMOVED_REG_7            (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKTS_REMOVED})
 `define OQ_ADDRESS_HI_REG_7                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_ADDRESS_HI})
 `define OQ_ADDRESS_LO_REG_7                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_ADDRESS_LO})
 `define OQ_WR_ADDRESS_REG_7                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_WR_ADDRESS})
 `define OQ_RD_ADDRESS_REG_7                  (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_RD_ADDRESS})
 `define OQ_NUM_PKTS_IN_Q_REG_7               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_PKTS_IN_Q})
 `define OQ_MAX_PKTS_IN_Q_REG_7               (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_MAX_PKTS_IN_Q})
 `define OQ_CONTROL_REG_7                     (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_CONTROL})
 `define OQ_FULL_THRESH_REG_7                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_FULL_THRESH})
 `define OQ_NUM_WORDS_IN_Q_REG_7              (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h7}, `OQ_NUM_WORDS_IN_Q})
 //////////////////////////////////////////////////
 `define JAN_OQ_BLOCK_CNT_REG7                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_BLOCK_CNT}) 
 `define JAN_OQ_PKTRM_CNT_REG7                (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_PKTRM_CNT})
 `define JAN_OQ_AB_STATE_REG7                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_STATE})
 `define JAN_OQ_AB_MOD_STATE_REG7             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AB_MOD_STATE})
 `define JAN_OQ_AC_STATE_REG7                 (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_STATE})
 `define JAN_OQ_AC_MOD_STATE_REG7             (`UDP_BASE_ADDRESS | {`OQ_BLOCK_TAG, {`OQ_REG_HELPER_BLOCK_ADDR_WIDTH'h0}, `JAN_OQ_AC_MOD_STATE})
//////////////////////////////////////////////////////////////////////////////////////////

 `define DELAY_ENABLE_REG                     (`UDP_BASE_ADDRESS | {`DELAY_BLOCK_TAG, `DELAY_ENABLE})
 `define DELAY_LENGTH_REG                     (`UDP_BASE_ADDRESS | {`DELAY_BLOCK_TAG, `DELAY_LENGTH})
 `define DELAY_1ST_WORD_HI_REG                (`UDP_BASE_ADDRESS | {`DELAY_BLOCK_TAG, `DELAY_1ST_WORD_HI})
 `define DELAY_1ST_WORD_LO_REG                (`UDP_BASE_ADDRESS | {`DELAY_BLOCK_TAG, `DELAY_1ST_WORD_LO})

 `define RATE_LIMIT_ENABLE_REG                (`UDP_BASE_ADDRESS | {`RATE_LIMIT_BLOCK_TAG, `RATE_LIMIT_ENABLE})
 `define RATE_LIMIT_SHIFT_REG                 (`UDP_BASE_ADDRESS | {`RATE_LIMIT_BLOCK_TAG, `RATE_LIMIT_SHIFT})

 `define EVT_CAP_ENABLE_CAPTURE_REG           (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_ENABLE_CAPTURE})
 `define EVT_CAP_SEND_PKT_REG                 (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_SEND_PKT})
 `define EVT_CAP_DST_MAC_HI_REG               (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_DST_MAC_HI})
 `define EVT_CAP_DST_MAC_LO_REG               (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_DST_MAC_LO})
 `define EVT_CAP_SRC_MAC_HI_REG               (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_SRC_MAC_HI})
 `define EVT_CAP_SRC_MAC_LO_REG               (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_SRC_MAC_LO})
 `define EVT_CAP_ETHERTYPE_REG                (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_ETHERTYPE})
 `define EVT_CAP_IP_DST_REG                   (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_IP_DST})
 `define EVT_CAP_IP_SRC_REG                   (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_IP_SRC})
 `define EVT_CAP_UDP_SRC_PORT_REG             (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_UDP_SRC_PORT})
 `define EVT_CAP_UDP_DST_PORT_REG             (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_UDP_DST_PORT})
 `define EVT_CAP_OUTPUT_PORTS_REG             (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_OUTPUT_PORTS})
 `define EVT_CAP_RESET_TIMERS_REG             (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_RESET_TIMERS})
 `define EVT_CAP_MONITOR_MASK_REG             (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_MONITOR_MASK})
 `define EVT_CAP_TIMER_RESOLUTION_REG         (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_TIMER_RESOLUTION})
 `define EVT_CAP_NUM_EVT_PKTS_SENT_REG        (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_NUM_EVT_PKTS_SENT})
 `define EVT_CAP_NUM_EVTS_SENT_REG            (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_NUM_EVTS_SENT})
 `define EVT_CAP_NUM_EVTS_DROPPED_REG         (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_NUM_EVTS_DROPPED})
 `define EVT_CAP_SIGNAL_ID_MASK_REG           (`UDP_BASE_ADDRESS | {`EVT_CAP_BLOCK_TAG, `EVT_CAP_SIGNAL_ID_MASK})

 `define DECAP_NUM_WORD_IN_REG                (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_NUM_WORD_IN})
 `define DECAP_NUM_WORD_OUT_REG               (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_NUM_WORD_OUT})
 `define DECAP_VALID_TUNNELING_REG            (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_VALID_TUNNELING})
 `define DECAP_USER_DATA_PATH_HEADER_REG      (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_USER_DATA_PATH_HEADER})
 `define DECAP_NUM_PACKET_IN_REG              (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_NUM_PACKET_IN})
 `define DECAP_NUM_PACKET_OUT_REG             (`UDP_BASE_ADDRESS | {`DECAP_BLOCK_TAG, `DECAP_NUM_PACKET_OUT})


 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_0_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_0})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_0_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_0})
 `define BRAM_OQ_NUM_PKTS_DROPPED_0_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_0})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_1_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_1})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_1_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_1})
 `define BRAM_OQ_NUM_PKTS_DROPPED_1_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_1})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_2_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_2})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_2_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_2})
 `define BRAM_OQ_NUM_PKTS_DROPPED_2_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_2})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_3_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_3})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_3_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_3})
 `define BRAM_OQ_NUM_PKTS_DROPPED_3_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_3})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_4_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_4})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_4_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_4})
 `define BRAM_OQ_NUM_PKTS_DROPPED_4_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_4})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_5_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_5})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_5_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_5})
 `define BRAM_OQ_NUM_PKTS_DROPPED_5_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_5})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_6_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_6})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_6_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_6})
 `define BRAM_OQ_NUM_PKTS_DROPPED_6_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_6})
 `define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_7_REG (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_7})
 `define BRAM_OQ_NUM_PKTS_RECEIVED_7_REG      (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_RECEIVED_7})
 `define BRAM_OQ_NUM_PKTS_DROPPED_7_REG       (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_PKTS_DROPPED_7})
 `define BRAM_OQ_DISABLE_QUEUES_REG           (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_DISABLE_QUEUES})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_0_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_0})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_1_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_1})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_2_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_2})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_3_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_3})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_4_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_4})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_5_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_5})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_6_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_6})
 `define BRAM_OQ_NUM_WORDS_IN_QUEUE_7_REG     (`UDP_BASE_ADDRESS | {`BRAM_OQ_BLOCK_TAG, `BRAM_OQ_NUM_WORDS_IN_QUEUE_7})
 
 `define RCP_RATE_REG                         (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_RATE})
 `define RCP_MAC_0_RTT_L_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_0_RTT_L})
 `define RCP_MAC_0_RTT_H_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_0_RTT_H})
 `define RCP_MAC_0_NUM_BYTE_L_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_0_NUM_BYTE_L})
 `define RCP_MAC_0_NUM_BYTE_H_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_0_NUM_BYTE_H})
 `define RCP_MAC_0_NUM_RCP_REG                (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_0_NUM_RCP})
 `define RCP_MAC_1_RTT_L_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_1_RTT_L})
 `define RCP_MAC_1_RTT_H_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_1_RTT_H})
 `define RCP_MAC_1_NUM_BYTE_L_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_1_NUM_BYTE_L})
 `define RCP_MAC_1_NUM_BYTE_H_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_1_NUM_BYTE_H})
 `define RCP_MAC_1_NUM_RCP_REG                (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_1_NUM_RCP})
 `define RCP_MAC_2_RTT_L_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_2_RTT_L})
 `define RCP_MAC_2_RTT_H_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_2_RTT_H})
 `define RCP_MAC_2_NUM_BYTE_L_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_2_NUM_BYTE_L})
 `define RCP_MAC_2_NUM_BYTE_H_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_2_NUM_BYTE_H})
 `define RCP_MAC_2_NUM_RCP_REG                (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_2_NUM_RCP})

 `define RCP_MAC_3_RTT_L_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_3_RTT_L})
 `define RCP_MAC_3_RTT_H_REG                  (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_3_RTT_H})
 `define RCP_MAC_3_NUM_BYTE_L_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_3_NUM_BYTE_L})
 `define RCP_MAC_3_NUM_BYTE_H_REG             (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_3_NUM_BYTE_H})
 `define RCP_MAC_3_NUM_RCP_REG                (`UDP_BASE_ADDRESS | {`RCP_BLOCK_TAG, `RCP_MAC_3_NUM_RCP})

 `define PKT_GEN_CTRL_ENABLE_REG              (`UDP_BASE_ADDRESS | {`PKT_GEN_CTRL_BLOCK_TAG, `PKT_GEN_CTRL_ENABLE})

 // 4- add external addresses here

 // ENCAP
 `define ENCAP_ENABLE_REG                      (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_ENABLE})
 `define ENCAP_IP_DATA_0_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_0})
 `define ENCAP_IP_DATA_1_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_1})
 `define ENCAP_IP_DATA_2_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_2})
 `define ENCAP_IP_DATA_3_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_3})
 `define ENCAP_IP_DATA_4_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_4})
 `define ENCAP_IP_DATA_5_REG                   (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_IP_DATA_5})
 `define ENCAP_NUM_PACKET_IN_REG               (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_NUM_PACKET_IN})
 `define ENCAP_NUM_PACKET_OUT_REG              (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_NUM_PACKET_OUT})
 `define ENCAP_NUM_BYTES_IN_REG                (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_NUM_BYTES_IN})
 `define ENCAP_NUM_BYTES_OUT_REG               (`UDP_BASE_ADDRESS  | {`ENCAP_BLOCK_TAG, `ENCAP_NUM_BYTES_OUT})


 /*********************************************************
 * useful macros
 *********************************************************/

 // 5- print the reg name and addr in C format
 `define PRINT_REG_ADDRESSES_UDP                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_NUM_PKTS_SENT_REG                  0x%07x\n", `IN_ARB_NUM_PKTS_SENT_REG<<2);                    \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_WORD_0_LO_REG             0x%07x\n", `IN_ARB_LAST_PKT_WORD_0_LO_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_WORD_0_HI_REG             0x%07x\n", `IN_ARB_LAST_PKT_WORD_0_HI_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_CTRL_0_REG                0x%07x\n", `IN_ARB_LAST_PKT_CTRL_0_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_WORD_1_LO_REG             0x%07x\n", `IN_ARB_LAST_PKT_WORD_1_LO_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_WORD_1_HI_REG             0x%07x\n", `IN_ARB_LAST_PKT_WORD_1_HI_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_LAST_PKT_CTRL_1_REG                0x%07x\n", `IN_ARB_LAST_PKT_CTRL_1_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define IN_ARB_STATE_REG                          0x%07x\n\n", `IN_ARB_STATE_REG<<2);                          \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_PORTS_MAC_HI_REG            0x%07x\n", `SWITCH_OP_LUT_PORTS_MAC_HI_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_MAC_LO_REG                  0x%07x\n", `SWITCH_OP_LUT_MAC_LO_REG<<2);                    \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_NUM_HITS_REG                0x%07x\n", `SWITCH_OP_LUT_NUM_HITS_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_NUM_MISSES_REG              0x%07x\n", `SWITCH_OP_LUT_NUM_MISSES_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_MAC_LUT_RD_ADDR_REG         0x%07x\n", `SWITCH_OP_LUT_MAC_LUT_RD_ADDR_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define SWITCH_OP_LUT_MAC_LUT_WR_ADDR_REG         0x%07x\n\n", `SWITCH_OP_LUT_MAC_LUT_WR_ADDR_REG<<2);         \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define ROUTER_RT_SIZE                            %d\n", `ROUTER_RT_SIZE);                                     \
         $fwrite(c_reg_defines_fd, "#define ROUTER_ARP_SIZE                           %d\n", `ROUTER_ARP_SIZE);                                    \
         $fwrite(c_reg_defines_fd, "#define ROUTER_DST_IP_FILTER_TABLE_DEPTH          %d\n\n", `ROUTER_DST_IP_FILTER_TABLE_DEPTH);                 \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_MAC_HI_REG              0x%07x\n", `ROUTER_OP_LUT_ARP_MAC_HI_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_MAC_LO_REG              0x%07x\n", `ROUTER_OP_LUT_ARP_MAC_LO_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_NEXT_HOP_IP_REG         0x%07x\n", `ROUTER_OP_LUT_ARP_NEXT_HOP_IP_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_LUT_RD_ADDR_REG         0x%07x\n", `ROUTER_OP_LUT_ARP_LUT_RD_ADDR_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_LUT_WR_ADDR_REG         0x%07x\n", `ROUTER_OP_LUT_ARP_LUT_WR_ADDR_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_IP_REG                   0x%07x\n", `ROUTER_OP_LUT_RT_IP_REG<<2);                     \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_MASK_REG                 0x%07x\n", `ROUTER_OP_LUT_RT_MASK_REG<<2);                   \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_NEXT_HOP_IP_REG          0x%07x\n", `ROUTER_OP_LUT_RT_NEXT_HOP_IP_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_OUTPUT_PORT_REG          0x%07x\n", `ROUTER_OP_LUT_RT_OUTPUT_PORT_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_LUT_RD_ADDR_REG          0x%07x\n", `ROUTER_OP_LUT_RT_LUT_RD_ADDR_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_RT_LUT_WR_ADDR_REG          0x%07x\n", `ROUTER_OP_LUT_RT_LUT_WR_ADDR_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_0_HI_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_0_HI_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_0_LO_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_0_LO_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_1_HI_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_1_HI_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_1_LO_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_1_LO_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_2_HI_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_2_HI_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_2_LO_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_2_LO_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_3_HI_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_3_HI_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_MAC_3_LO_REG                0x%07x\n", `ROUTER_OP_LUT_MAC_3_LO_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_DST_IP_FILTER_IP_REG        0x%07x\n", `ROUTER_OP_LUT_DST_IP_FILTER_IP_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_DST_IP_FILTER_RD_ADDR_REG   0x%07x\n", `ROUTER_OP_LUT_DST_IP_FILTER_RD_ADDR_REG<<2);     \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_DST_IP_FILTER_WR_ADDR_REG   0x%07x\n\n", `ROUTER_OP_LUT_DST_IP_FILTER_WR_ADDR_REG<<2);   \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_ARP_NUM_MISSES_REG          0x%07x\n", `ROUTER_OP_LUT_ARP_NUM_MISSES_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_LPM_NUM_MISSES_REG          0x%07x\n", `ROUTER_OP_LUT_LPM_NUM_MISSES_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_CPU_PKTS_SENT_REG       0x%07x\n", `ROUTER_OP_LUT_NUM_CPU_PKTS_SENT_REG<<2);         \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_BAD_OPTS_VER_REG        0x%07x\n", `ROUTER_OP_LUT_NUM_BAD_OPTS_VER_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_BAD_CHKSUMS_REG         0x%07x\n", `ROUTER_OP_LUT_NUM_BAD_CHKSUMS_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_BAD_TTLS_REG            0x%07x\n", `ROUTER_OP_LUT_NUM_BAD_TTLS_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_NON_IP_RCVD_REG         0x%07x\n", `ROUTER_OP_LUT_NUM_NON_IP_RCVD_REG<<2);           \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_PKTS_FORWARDED_REG      0x%07x\n", `ROUTER_OP_LUT_NUM_PKTS_FORWARDED_REG<<2);        \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_WRONG_DEST_REG          0x%07x\n", `ROUTER_OP_LUT_NUM_WRONG_DEST_REG<<2);            \
         $fwrite(c_reg_defines_fd, "#define ROUTER_OP_LUT_NUM_FILTERED_PKTS_REG       0x%07x\n\n", `ROUTER_OP_LUT_NUM_FILTERED_PKTS_REG<<2);       \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define OQ_ENABLE_SEND_BIT_NUM                    %d\n", `OQ_ENABLE_SEND_BIT_NUM);                             \
         $fwrite(c_reg_defines_fd, "#define OQ_INITIALIZE_OQ_BIT_NUM                  %d\n\n", `OQ_INITIALIZE_OQ_BIT_NUM);                         \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_0                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_0<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_0           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_0<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_0      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_0<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_0                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_0<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_0               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_0<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_0          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_0<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_0     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_0<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_0               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_0<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_0                     0x%07x\n", `OQ_ADDRESS_HI_REG_0<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_0                     0x%07x\n", `OQ_ADDRESS_LO_REG_0<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_0                     0x%07x\n", `OQ_WR_ADDRESS_REG_0<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_0                     0x%07x\n", `OQ_RD_ADDRESS_REG_0<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_0                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_0<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_0                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_0<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_0                    0x%07x\n", `OQ_FULL_THRESH_REG_0<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_0                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_0<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_0                        0x%07x\n\n", `OQ_CONTROL_REG_0<<2);                            \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG0                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG0<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG0                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG0<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG0                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG0<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG0                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG0<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG0                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG0<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG0                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG0<<2);                    \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_1                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_1<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_1           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_1<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_1      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_1<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_1                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_1<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_1               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_1<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_1          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_1<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_1     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_1<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_1               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_1<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_1                     0x%07x\n", `OQ_ADDRESS_HI_REG_1<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_1                     0x%07x\n", `OQ_ADDRESS_LO_REG_1<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_1                     0x%07x\n", `OQ_WR_ADDRESS_REG_1<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_1                     0x%07x\n", `OQ_RD_ADDRESS_REG_1<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_1                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_1<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_1                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_1<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_1                    0x%07x\n", `OQ_FULL_THRESH_REG_1<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_1                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_1<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_1                        0x%07x\n\n", `OQ_CONTROL_REG_1<<2);                            \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG1                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG1<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG1                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG1<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG1                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG1<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG1                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG1<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG1                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG1<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG1                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG1<<2);                    \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_2                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_2<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_2           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_2<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_2      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_2<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_2                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_2<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_2               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_2<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_2          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_2<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_2     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_2<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_2               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_2<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_2                     0x%07x\n", `OQ_ADDRESS_HI_REG_2<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_2                     0x%07x\n", `OQ_ADDRESS_LO_REG_2<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_2                     0x%07x\n", `OQ_WR_ADDRESS_REG_2<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_2                     0x%07x\n", `OQ_RD_ADDRESS_REG_2<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_2                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_2<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_2                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_2<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_2                    0x%07x\n", `OQ_FULL_THRESH_REG_2<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_2                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_2<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_2                        0x%07x\n\n", `OQ_CONTROL_REG_2<<2);                            \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG2                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG2<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG2                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG2<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG2                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG2<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG2                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG2<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG2                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG2<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG2                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG2<<2);                    \		                                                                                                                                                    \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_3                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_3<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_3           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_3<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_3      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_3<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_3                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_3<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_3               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_3<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_3          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_3<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_3     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_3<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_3               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_3<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_3                     0x%07x\n", `OQ_ADDRESS_HI_REG_3<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_3                     0x%07x\n", `OQ_ADDRESS_LO_REG_3<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_3                     0x%07x\n", `OQ_WR_ADDRESS_REG_3<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_3                     0x%07x\n", `OQ_RD_ADDRESS_REG_3<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_3                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_3<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_3                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_3<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_3                    0x%07x\n", `OQ_FULL_THRESH_REG_3<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_3                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_3<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_3                        0x%07x\n\n", `OQ_CONTROL_REG_3<<2);                            \
		 $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG3                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG3<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG3                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG3<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG3                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG3<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG3                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG3<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG3                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG3<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG3                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG3<<2);                    \                                                                                                                                                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_4                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_4<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_4           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_4<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_4      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_4<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_4                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_4<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_4               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_4<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_4          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_4<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_4     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_4<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_4               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_4<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_4                     0x%07x\n", `OQ_ADDRESS_HI_REG_4<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_4                     0x%07x\n", `OQ_ADDRESS_LO_REG_4<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_4                     0x%07x\n", `OQ_WR_ADDRESS_REG_4<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_4                     0x%07x\n", `OQ_RD_ADDRESS_REG_4<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_4                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_4<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_4                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_4<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_4                    0x%07x\n", `OQ_FULL_THRESH_REG_4<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_4                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_4<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_4                        0x%07x\n\n", `OQ_CONTROL_REG_4<<2);                            \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG4                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG4<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG4                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG4<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG4                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG4<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG4                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG4<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG4                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG4<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG4                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG4<<2);                    \
	  	                                                                                                                                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_5                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_5<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_5           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_5<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_5      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_5<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_5                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_5<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_5               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_5<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_5          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_5<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_5     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_5<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_5               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_5<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_5                     0x%07x\n", `OQ_ADDRESS_HI_REG_5<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_5                     0x%07x\n", `OQ_ADDRESS_LO_REG_5<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_5                     0x%07x\n", `OQ_WR_ADDRESS_REG_5<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_5                     0x%07x\n", `OQ_RD_ADDRESS_REG_5<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_5                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_5<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_5                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_5<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_5                    0x%07x\n", `OQ_FULL_THRESH_REG_5<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_5                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_5<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_5                        0x%07x\n\n", `OQ_CONTROL_REG_5<<2);                            \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG5                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG5<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG5                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG5<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG5                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG5<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG5                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG5<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG5                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG5<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG5                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG5<<2);                    \
                                                                                                                                            	  \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_6                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_6<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_6           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_6<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_6      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_6<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_6                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_6<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_6               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_6<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_6          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_6<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_6     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_6<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_6               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_6<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_6                     0x%07x\n", `OQ_ADDRESS_HI_REG_6<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_6                     0x%07x\n", `OQ_ADDRESS_LO_REG_6<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_6                     0x%07x\n", `OQ_WR_ADDRESS_REG_6<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_6                     0x%07x\n", `OQ_RD_ADDRESS_REG_6<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_6                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_6<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_6                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_6<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_6                    0x%07x\n", `OQ_FULL_THRESH_REG_6<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_6                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_6<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_6                        0x%07x\n\n", `OQ_CONTROL_REG_6<<2);                            \
		 $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG6                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG6<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG6                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG6<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG6                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG6<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG6                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG6<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG6                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG6<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG6                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG6<<2);                    \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_LEFT_REG_7                 0x%07x\n", `OQ_NUM_WORDS_LEFT_REG_7<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_STORED_REG_7           0x%07x\n", `OQ_NUM_PKT_BYTES_STORED_REG_7<<2);                 \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_STORED_REG_7      0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_STORED_REG_7<<2);            \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_STORED_REG_7                0x%07x\n", `OQ_NUM_PKTS_STORED_REG_7<<2);                      \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_DROPPED_REG_7               0x%07x\n", `OQ_NUM_PKTS_DROPPED_REG_7<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKT_BYTES_REMOVED_REG_7          0x%07x\n", `OQ_NUM_PKT_BYTES_REMOVED_REG_7<<2);                \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_7     0x%07x\n", `OQ_NUM_OVERHEAD_BYTES_REMOVED_REG_7<<2);           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_REMOVED_REG_7               0x%07x\n", `OQ_NUM_PKTS_REMOVED_REG_7<<2);                     \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_HI_REG_7                     0x%07x\n", `OQ_ADDRESS_HI_REG_7<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_ADDRESS_LO_REG_7                     0x%07x\n", `OQ_ADDRESS_LO_REG_7<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_WR_ADDRESS_REG_7                     0x%07x\n", `OQ_WR_ADDRESS_REG_7<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_RD_ADDRESS_REG_7                     0x%07x\n", `OQ_RD_ADDRESS_REG_7<<2);                           \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_PKTS_IN_Q_REG_7                  0x%07x\n", `OQ_NUM_PKTS_IN_Q_REG_7<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_MAX_PKTS_IN_Q_REG_7                  0x%07x\n", `OQ_MAX_PKTS_IN_Q_REG_7<<2);                        \
         $fwrite(c_reg_defines_fd, "#define OQ_FULL_THRESH_REG_7                    0x%07x\n", `OQ_FULL_THRESH_REG_7<<2);                          \
         $fwrite(c_reg_defines_fd, "#define OQ_NUM_WORDS_IN_Q_REG_7                 0x%07x\n", `OQ_NUM_WORDS_IN_Q_REG_7<<2);                       \
         $fwrite(c_reg_defines_fd, "#define OQ_CONTROL_REG_7                        0x%07x\n\n", `OQ_CONTROL_REG_7<<2);                            \
		 $fwrite(c_reg_defines_fd, "#define JAN_OQ_BLOCK_CNT_REG7                   0x%07x\n\n", `JAN_OQ_BLOCK_CNT_REG7<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_PKTRM_CNT_REG7                   0x%07x\n\n", `JAN_OQ_PKTRM_CNT_REG7<<2);                       \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_STATE_REG7                    0x%07x\n\n", `JAN_OQ_AB_STATE_REG7<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AB_MOD_STATE_REG7                0x%07x\n\n", `JAN_OQ_AB_MOD_STATE_REG7<<2);                    \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_STATE_REG7                    0x%07x\n\n", `JAN_OQ_AC_STATE_REG7<<2);                        \
         $fwrite(c_reg_defines_fd, "#define JAN_OQ_AC_MOD_STATE_REG7                0x%07x\n\n", `JAN_OQ_AC_MOD_STATE_REG7<<2);                    \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define DELAY_ENABLE_REG                        0x%07x\n", `DELAY_ENABLE_REG<<2);                              \
         $fwrite(c_reg_defines_fd, "#define DELAY_1ST_WORD_HI_REG                   0x%07x\n", `DELAY_1ST_WORD_HI_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define DELAY_1ST_WORD_LO_REG                   0x%07x\n", `DELAY_1ST_WORD_LO_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define DELAY_LENGTH_REG                        0x%07x\n\n", `DELAY_LENGTH_REG<<2);                            \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define RATE_LIMIT_ENABLE_REG                   0x%07x\n", `RATE_LIMIT_ENABLE_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define RATE_LIMIT_SHIFT_REG                    0x%07x\n\n", `RATE_LIMIT_SHIFT_REG<<2);                        \
                                                                                                                                                   \
         $fwrite(c_reg_defines_fd, "#define RCP_RATE_REG                            0x%07x\n", `RCP_RATE_REG<<2);                                  \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_0_RTT_L_REG                     0x%07x\n", `RCP_MAC_0_RTT_L_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_0_RTT_H_REG                     0x%07x\n", `RCP_MAC_0_RTT_H_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_0_NUM_RCP_REG                   0x%07x\n", `RCP_MAC_0_NUM_RCP_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_0_NUM_BYTE_L_REG                0x%07x\n", `RCP_MAC_0_NUM_BYTE_L_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_0_NUM_BYTE_H_REG                0x%07x\n", `RCP_MAC_0_NUM_BYTE_H_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_1_RTT_L_REG                     0x%07x\n", `RCP_MAC_1_RTT_L_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_1_RTT_H_REG                     0x%07x\n", `RCP_MAC_1_RTT_H_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_1_NUM_RCP_REG                   0x%07x\n", `RCP_MAC_1_NUM_RCP_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_1_NUM_BYTE_L_REG                0x%07x\n", `RCP_MAC_1_NUM_BYTE_L_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_1_NUM_BYTE_H_REG                0x%07x\n", `RCP_MAC_1_NUM_BYTE_H_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_2_RTT_L_REG                     0x%07x\n", `RCP_MAC_2_RTT_L_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_2_RTT_H_REG                     0x%07x\n", `RCP_MAC_2_RTT_H_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_2_NUM_RCP_REG                   0x%07x\n", `RCP_MAC_2_NUM_RCP_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_2_NUM_BYTE_L_REG                0x%07x\n", `RCP_MAC_2_NUM_BYTE_L_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_2_NUM_BYTE_H_REG                0x%07x\n", `RCP_MAC_2_NUM_BYTE_H_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_3_RTT_L_REG                     0x%07x\n", `RCP_MAC_3_RTT_L_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_3_RTT_H_REG                     0x%07x\n", `RCP_MAC_3_RTT_H_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_3_NUM_RCP_REG                   0x%07x\n\n", `RCP_MAC_3_NUM_RCP_REG<<2);                       \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_3_NUM_BYTE_L_REG                0x%07x\n", `RCP_MAC_3_NUM_BYTE_L_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define RCP_MAC_3_NUM_BYTE_H_REG                0x%07x\n", `RCP_MAC_3_NUM_BYTE_H_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_ENABLE_CAPTURE_REG              0x%07x\n", `EVT_CAP_ENABLE_CAPTURE_REG<<2);                    \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_SEND_PKT_REG                    0x%07x\n", `EVT_CAP_SEND_PKT_REG<<2);                          \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_DST_MAC_HI_REG                  0x%07x\n", `EVT_CAP_DST_MAC_HI_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_DST_MAC_LO_REG                  0x%07x\n", `EVT_CAP_DST_MAC_LO_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_SRC_MAC_HI_REG                  0x%07x\n", `EVT_CAP_SRC_MAC_HI_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_SRC_MAC_LO_REG                  0x%07x\n", `EVT_CAP_SRC_MAC_LO_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_ETHERTYPE_REG                   0x%07x\n", `EVT_CAP_ETHERTYPE_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_IP_DST_REG                      0x%07x\n", `EVT_CAP_IP_DST_REG<<2);                            \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_IP_SRC_REG                      0x%07x\n", `EVT_CAP_IP_SRC_REG<<2);                            \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_UDP_SRC_PORT_REG                0x%07x\n", `EVT_CAP_UDP_SRC_PORT_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_UDP_DST_PORT_REG                0x%07x\n", `EVT_CAP_UDP_DST_PORT_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_OUTPUT_PORTS_REG                0x%07x\n", `EVT_CAP_OUTPUT_PORTS_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_RESET_TIMERS_REG                0x%07x\n", `EVT_CAP_RESET_TIMERS_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_MONITOR_MASK_REG                0x%07x\n", `EVT_CAP_MONITOR_MASK_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_TIMER_RESOLUTION_REG            0x%07x\n", `EVT_CAP_TIMER_RESOLUTION_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_NUM_EVT_PKTS_SENT_REG           0x%07x\n", `EVT_CAP_NUM_EVT_PKTS_SENT_REG<<2);                 \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_NUM_EVTS_SENT_REG               0x%07x\n", `EVT_CAP_NUM_EVTS_SENT_REG<<2);                     \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_NUM_EVTS_DROPPED_REG            0x%07x\n", `EVT_CAP_NUM_EVTS_DROPPED_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define EVT_CAP_SIGNAL_ID_MASK_REG              0x%07x\n\n", `EVT_CAP_SIGNAL_ID_MASK_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define DECAP_NUM_WORD_IN_REG                   0x%07x\n", `DECAP_NUM_WORD_IN_REG<<2);                         \
         $fwrite(c_reg_defines_fd, "#define DECAP_NUM_WORD_OUT_REG                  0x%07x\n", `DECAP_NUM_WORD_OUT_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define DECAP_VALID_TUNNELING_REG               0x%07x\n", `DECAP_VALID_TUNNELING_REG<<2);                     \
         $fwrite(c_reg_defines_fd, "#define DECAP_USER_DATA_PATH_HEADER_REG         0x%07x\n", `DECAP_USER_DATA_PATH_HEADER_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define DECAP_NUM_PACKET_IN_REG                 0x%07x\n", `DECAP_NUM_PACKET_IN_REG<<2);                       \
         $fwrite(c_reg_defines_fd, "#define DECAP_NUM_PACKET_OUT_REG                0x%07x\n", `DECAP_NUM_PACKET_OUT_REG<<2);                      \
         $fwrite(c_reg_defines_fd, "#define ENCAP_NUM_PACKET_IN_REG                   0x%07x\n\n", `ENCAP_NUM_PACKET_IN_REG<<2);                   \
	$fwrite(c_reg_defines_fd, "#define ENCAP_NUM_PACKET_OUT_REG                   0x%07x\n\n", `ENCAP_NUM_PACKET_OUT_REG<<2);                  \
         $fwrite(c_reg_defines_fd, "#define ENCAP_NUM_BYTES_IN_REG                 0x%07x\n\n", `ENCAP_NUM_BYTES_IN_REG<<2);                       \
         $fwrite(c_reg_defines_fd, "#define ENCAP_NUM_BYTES_OUT_REG                 0x%07x\n\n", `ENCAP_NUM_BYTES_OUT_REG<<2);                    \
	 $fwrite(c_reg_defines_fd, "#define ENCAP_ENABLE_REG                        0x%07x\n\n", `ENCAP_ENABLE_REG<<2);                           \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_0_REG                     0x%07x\n\n", `ENCAP_IP_DATA_0_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_1_REG                     0x%07x\n\n", `ENCAP_IP_DATA_1_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_2_REG                     0x%07x\n\n", `ENCAP_IP_DATA_2_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_3_REG                     0x%07x\n\n", `ENCAP_IP_DATA_3_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_4_REG                     0x%07x\n\n", `ENCAP_IP_DATA_4_REG<<2);                        \
         $fwrite(c_reg_defines_fd, "#define ENCAP_IP_DATA_5_REG                     0x%07x\n\n", `ENCAP_IP_DATA_5_REG<<2);                        \
        $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_0_REG     0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_0_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_0_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_0_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_0_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_0_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_1_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_1_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_1_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_1_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_1_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_1_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_2_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_2_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_2_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_2_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_2_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_2_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_3_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_3_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_3_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_3_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_3_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_3_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_4_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_4_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_4_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_4_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_4_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_4_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_5_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_5_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_5_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_5_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_5_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_5_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_6_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_6_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_6_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_6_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_6_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_6_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKT_BYTES_RECEIVED_7_REG    0x%07x\n", `BRAM_OQ_NUM_PKT_BYTES_RECEIVED_7_REG<<2);          \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_RECEIVED_7_REG         0x%07x\n", `BRAM_OQ_NUM_PKTS_RECEIVED_7_REG<<2);               \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_PKTS_DROPPED_7_REG          0x%07x\n", `BRAM_OQ_NUM_PKTS_DROPPED_7_REG<<2);                \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_DISABLE_QUEUES_REG              0x%07x\n", `BRAM_OQ_DISABLE_QUEUES_REG<<2);                    \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_0_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_0_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_1_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_1_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_2_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_2_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_3_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_3_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_4_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_4_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_5_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_5_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_6_REG        0x%07x\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_6_REG<<2);              \
         $fwrite(c_reg_defines_fd, "#define BRAM_OQ_NUM_WORDS_IN_QUEUE_7_REG        0x%07x\n\n", `BRAM_OQ_NUM_WORDS_IN_QUEUE_7_REG<<2)
                                                              
`endif //  `ifndef _UDP_DEFINES_


