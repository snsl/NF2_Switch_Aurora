//
//      Project:  Aurora Module Generator version 2.9
//
//         Date:  $Date: 2007/10/04 04:15:13 $
//          Tag:  $Name: i+IP+138572 $
//         File:  $RCSfile: frame_check.ejava,v $
//          Rev:  $Revision: 1.1.2.1 $
//
//      Company:  Xilinx
//
//   Disclaimer:  XILINX IS PROVIDING THIS DESIGN, CODE, OR
//                INFORMATION "AS IS" SOLELY FOR USE IN DEVELOPING
//                PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY
//                PROVIDING THIS DESIGN, CODE, OR INFORMATION AS
//                ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE,
//                APPLICATION OR STANDARD, XILINX IS MAKING NO
//                REPRESENTATION THAT THIS IMPLEMENTATION IS FREE
//                FROM ANY CLAIMS OF INFRINGEMENT, AND YOU ARE
//                RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY
//                REQUIRE FOR YOUR IMPLEMENTATION.  XILINX
//                EXPRESSLY DISCLAIMS ANY WARRANTY WHATSOEVER WITH
//                RESPECT TO THE ADEQUACY OF THE IMPLEMENTATION,
//                INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR
//                REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE
//                FROM CLAIMS OF INFRINGEMENT, IMPLIED WARRANTIES
//                OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
//                PURPOSE.
//
//                (c) Copyright 2004 Xilinx, Inc.
//                All rights reserved.
//

//
//  FRAME CHECK
//
//
//
//  Description: This module is a  pattern checker to test the Aurora
//               designs in hardware. The frames generated by FRAME_GEN
//               pass through the Aurora channel and arrive at the frame checker 
//               through the RX User interface. Every time an error is found in
//               the data recieved, the error count is incremented until it 
//               reaches its max value.

`timescale 1 ns / 10 ps
`define DLY #1


module aurora_link_FRAME_CHECK
(
    // User Interface
    RX_D,  
    RX_REM,     
    RX_SOF_N,       
    RX_EOF_N,
    RX_SRC_RDY_N,  

    // System Interface
    USER_CLK,       
    RESET,
    ERROR_COUNT
  
);

//***********************************Port Declarations*******************************

   // User Interface
    input   [0:15]     RX_D;
    input              RX_REM;
    input              RX_SOF_N;
    input              RX_EOF_N;
    input              RX_SRC_RDY_N;
    
      // System Interface
    input              USER_CLK;
    input              RESET; 
    output  [0:7]      ERROR_COUNT;


//***************************Internal Register Declarations*************************** 

    reg                in_frame_r;
    reg     [0:15]     data_r;
    reg                data_valid_r;
    reg                error_detected_r;
    reg     [0:8]      error_count_r;
    
 
//*********************************Wire Declarations**********************************
   
    wire               data_valid_c;
    wire               in_frame_c;
    wire               rem_valid_c;
    
    wire               error_detected_c;


//*********************************Main Body of Code**********************************


    


    //______________________________ Capture incoming data ___________________________    
    //Data is valid when RX_SRC_RDY_N is asserted and data is arriving within a frame
    assign  data_valid_c    =   in_frame_c && rem_valid_c && !RX_SRC_RDY_N;


    //Data is in a frame if it is a single cycle frame or a multi_cycle frame has started
    assign  in_frame_c  =   in_frame_r  ||  (!RX_SRC_RDY_N && !RX_SOF_N);
    
    
    //Start a multicycle frame when a frame starts without ending on the same cycle. End 
    //the frame when an EOF is detected
    always @(posedge USER_CLK)
        if(RESET)   
            in_frame_r  <=  `DLY    1'b0;
        else if(!in_frame_r && !RX_SOF_N && !RX_SRC_RDY_N && RX_EOF_N)
            in_frame_r  <=  `DLY    1'b1;
        else if(in_frame_r && !RX_SRC_RDY_N && !RX_EOF_N)
            in_frame_r  <=  `DLY    1'b0;
            
            
    //We expect rem to indicate a full word of data on the EOF cycle
    assign  rem_valid_c =   RX_EOF_N || (RX_REM == 1'd1);
                


    //Capture valid incoming data, right shifted 1 bit for comparison with the next valid
    //incoming data
    always @(posedge USER_CLK)
        if(data_valid_c)    
            data_r  <=  `DLY    {RX_D[15],RX_D[0:14]};



    //Data in the data register is valid only if it was valid when captured and had no error
    always @(posedge USER_CLK)
        if(RESET)   data_valid_r    <=  `DLY    1'b0;
        else        data_valid_r    <=  `DLY    data_valid_c && !error_detected_c;



    
    //___________________________ Check incoming data for errors __________________________
         
    
    //An error is detected when valid data from the data register, when right shifted, does not match valid data
    //from the Aurora RX port
    assign  error_detected_c    =   data_valid_c && data_valid_r && (RX_D != data_r);   
    
    
    //We register the error_detected signal for use with the error counter logic
    always @(posedge USER_CLK)
        if(RESET)  
            error_detected_r    <=  `DLY    1'b0;
        else
            error_detected_r    <=  `DLY    error_detected_c;  

    
    
    //We count the total number of errors we detect. By keeping a count we make it less likely that we will miss
    //errors we did not directly observe. This counter must be reset when it reaches its max value
    always @(posedge USER_CLK)
        if(RESET)
            error_count_r       <=  `DLY    9'd0;
        else if(error_detected_r && !error_count_r[0] )
            error_count_r       <=  `DLY    error_count_r + 1;
            
    
    
    //Here we connect the lower 8 bits of the count (the MSbit is used only to check when the counter reaches
    //max value) to the module output
    assign  ERROR_COUNT =   error_count_r[1:8];
    
    
endmodule           
